*  Generated for: HSPICE
*  Design library name: takemura
*  Design cell name: sram
*  Design view name: sram
.option search='/home/takemura/Workspace/takemura'

.option MCBRIEF=2
.param vtn=AGAUSS(0.6,0,1.0) vtp=AGAUSS(0.6,0,1.0)
.option PARHIER = LOCAL
.include '/home/takemura/Workspace/takemura/addfile.txt'
.option ARTIST=2 PSF=2
.temp 25
.include 'modified02_45nm_bulk_BSIM4_v1.0_HSPICE_pm.txt'
*Custom Designer (TM) Version J-2014.12-SP2-2
*Mon Jul  2 16:21:08 2018

.GLOBAL gnd! vdd!
********************************************************************************
* Library          : takemura
* Cell             : sram
* View             : sram
* View Search List : hspice hspiceD schematic spice veriloga
* View Stop List   : hspice hspiceD
********************************************************************************
m30 m8d m7d vdd! vdd! PCH w=90n l=0.045u ad='(90n*0.14u)' as='(90n*0.14u)' pd='(2*(90n+0.14u))'
+  ps='(2*(90n+0.14u))'
m9 m7d m8d vdd! vdd! PCH w=90n l=0.045u ad='(90n*0.14u)' as='(90n*0.14u)' pd='(2*(90n+0.14u))'
+  ps='(2*(90n+0.14u))'
m31 blb v3 vdd! vdd! PCH1 w=90n l=0.045u ad='(90n*0.14u)' as='(90n*0.14u)' pd='(2*(90n+0.14u))'
+  ps='(2*(90n+0.14u))'
m32 bl v3 vdd! vdd! PCH1 w=90n l=0.045u ad='(90n*0.14u)' as='(90n*0.14u)' pd='(2*(90n+0.14u))'
+  ps='(2*(90n+0.14u))'
m27 m8d v2 bl gnd! NCH w=60n l=0.045u ad='(60n*0.14u)' as='(60n*0.14u)' pd='(2*(60n+0.14u))'
+  ps='(2*(60n+0.14u))'
m26 m8d m7d gnd! gnd! NCH w=60n l=0.045u ad='(60n*0.14u)' as='(60n*0.14u)' pd='(2*(60n+0.14u))'
+  ps='(2*(60n+0.14u))'
m24 bl v1 gnd! gnd! NCH1 w=300n l=0.045u ad='(300n*0.14u)' as='(300n*0.14u)' pd='(2*(300n+0.14u))'
+  ps='(2*(300n+0.14u))'
m14 blb gnd! gnd! gnd! NCH1 w=300n l=0.045u ad='(300n*0.14u)' as='(300n*0.14u)'
+ pd='(2*(300n+0.14u))' ps='(2*(300n+0.14u))'
m13 m7d v2 blb gnd! NCH w=60n l=0.045u ad='(60n*0.14u)' as='(60n*0.14u)' pd='(2*(60n+0.14u))'
+  ps='(2*(60n+0.14u))'
m25 m7d m8d gnd! gnd! NCH w=60n l=0.045u ad='(60n*0.14u)' as='(60n*0.14u)' pd='(2*(60n+0.14u))'
+  ps='(2*(60n+0.14u))'
v18 vdd! v1 dc=0 pulse ( 0.8 0 4.75n 0.5n 0.5n 9.5n 20n )
v35 vdd! v2 dc=0 pulse ( 0.8 0 4.75n 0.5n 0.5n 9.5n 20n )
v36 vdd! v3 dc=0 pulse ( 0.8 0 4.75n 0.5n 0.5n 9.5n 20n )





.tran 10p 20n start=0 uic sweep monte=100 firstrun=1
.option opfile=1 split_dp=2




.end